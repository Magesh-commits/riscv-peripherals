module i2c(
clk,
SCL,
SDA,
RST,
LEDG,
LEDR,
SW_1
);
input SCL,RST;//asynchronous reset input
input clk;
inout SDA;
input SW_1;
output [7:0] LEDG;
output [17:0] LEDR;
parameter [2:0] STATE_IDLE      = 3'h0,//idle
                STATE_DEV_ADDR  = 3'h1,//the slave addr match
                STATE_READ      = 3'h2,//the op=read 
                STATE_IDX_PTR   = 3'h3,//get the index of inner-register
                STATE_WRITE     = 3'h4;//write the data in the reg 


reg             start_detect;
reg             start_resetter;

reg             stop_detect;
reg             stop_resetter;

reg [3:0]       bit_counter;//(from 0 to 8)9counters-> one byte=8bits and one ack=1bit
reg [7:0]       input_shift;
reg             master_ack;
reg [2:0]       state;
reg [7:0]       reg_00,reg_01,reg_02;//slave_reg
reg [15:0]      conv,conf,lot,hit;
conv = 16'b0000000000000000;    //0000h
conf = 16'b1000010110000011;    //8583h
lot  = 16'b1000000000000000;    //8000h
hit  = 16'b0111111111111111;    //7fffh
localparam [11:0] i1 = 12'd3,
                  i2 = 12'd4,
                  i3 = 12'd5,
                  i4 = 12'd6,
                  i5 = 12'd7,
                  i6 = 12'd8,
                  i7 = 12'd9,
                  i8 = 12'd10;

reg [7:0]       output_shift;
reg             output_control;
reg [7:0]       index_pointer;
reg conv_loaded = 1'b0; 
always @(*) begin
    if (conv_loaded == 1) begin
        if (conv[15:4] < lot[15:4]) begin
            $display("ERROR: the input data is lower than the limit at time %0t", $time);
            $finish;
        end
        else if (conv[15:4] > hit[15:4]) begin
            $display("ERROR: the input data is higher than the limit at time %0t", $time);
            $finish;
        end
        else begin
            $display("Value within limits: %b", conv[15:4]);
        end
    end
end



parameter [6:0] device_address = 7'h48;
wire            start_rst = RST | start_resetter;//detect the START for one cycle
wire            stop_rst = RST | stop_resetter;//detect the STOP for one cycle
wire            lsb_bit = (bit_counter == 4'h7) && !start_detect;//the 8bits one byte data
wire            ack_bit = (bit_counter == 4'h8) && !start_detect;//the 9bites ack 
wire            address_detect = (input_shift[7:1] == device_address);//the input address match the slave
wire            read_write_bit = input_shift[0];// the write or read operation 0=write and 1=read
wire            write_strobe = (state == STATE_WRITE) && ack_bit;//write state and finish one byte=8bits
assign          SDA = output_control ? 1'bz : 1'b0;

//-----------------for LED------------------------
wire [7:0] LEDG;
wire [17:0] LEDR;

assign LEDG[7]=start_detect;
assign LEDG[6]=stop_detect;
assign LEDG[5]=1'b0;
assign LEDG[4]=master_ack;
assign LEDG[3]=1'b0;
assign LEDG[2:0]=state;

assign LEDR[17:14]=bit_counter;
assign LEDR[10]=SW_1;
assign LEDR[7:0]=reg_01;

//---------------------------------------------
//---------------detect the start--------------
//---------------------------------------------
always @ (posedge start_rst or negedge SDA)
begin
        if (start_rst)
                start_detect <= 1'b0;
        else
                start_detect <= SCL;
end

always @ (posedge RST or posedge SCL)
begin
        if (RST)
                start_resetter <= 1'b0;
        else
                start_resetter <= start_detect;
end
//the START just last for one cycle of SCL



//---------------------------------------------
//---------------detect the stop---------------
//---------------------------------------------
always @ (posedge stop_rst or posedge SDA)
begin   
        if (stop_rst)
                stop_detect <= 1'b0;
        else
                stop_detect <= SCL;
end

always @ (posedge RST or posedge SCL)
begin   
        if (RST)
                stop_resetter <= 1'b0;
        else
                stop_resetter <= stop_detect;
end
//the STOP just last for one cycle of SCL
//don't need to check the RESTART,due to: a START before it is STOP,it's START; 
//                                        a START before it is START,it's RESTART;
//the RESET and START combine can be recognise the RESTART,but it's doesn't matter



//---------------------------------------------
//---------------latch the data---------------
//---------------------------------------------
always @ (negedge SCL)
begin
        if (ack_bit || start_detect)
                bit_counter <= 4'h0;
        else
                bit_counter <= bit_counter + 4'h1;
end
//counter to 9(from 0 to 8), one byte=8bits and one ack 
always @ (posedge SCL)
        if (!ack_bit)
                input_shift <= {input_shift[6:0], SDA};
//at posedge SCL the data is stable,the input_shift get one byte=8bits



//---------------------------------------------
//------------slave-to-master transfer---------
//---------------------------------------------
always @ (posedge SCL)
        if (ack_bit)
                master_ack <= ~SDA;//the ack SDA is low
//the 9th bits= ack if the SDA=1'b0 it's a ACK, 



//---------------------------------------------
//------------state machine--------------------
//---------------------------------------------
always @ (posedge RST or negedge SCL)//jcyuan comment
begin
        if (RST)
                state <= STATE_IDLE;
        else if (start_detect)
                state <= STATE_DEV_ADDR;
        else if (ack_bit)//at the 9th cycle and change the state by ACK
        begin
                case (state)
                STATE_IDLE:
                        state <= STATE_IDLE;

                STATE_DEV_ADDR:
                        if (!address_detect)//addr don't match
                                state <= STATE_IDLE;
                        else if (read_write_bit)// addr match and operation is read
                                state <= STATE_READ;
                        else//addr match and operation is write
                                state <= STATE_IDX_PTR;

                STATE_READ:
                        if (master_ack)//get the master ack 
                                state <= STATE_READ;
                        else//no master ack ready to STOP
                                state <= STATE_IDLE;

                STATE_IDX_PTR:
                        state <= STATE_WRITE;//get the index and ready to write 

                STATE_WRITE:
                        state <= STATE_WRITE;//when the state is write the state 
                endcase
        end
        //if don't write and master send a stop,need to jump idle
        //the stop_detect is the next cycle of ACK
        else if(stop_detect)//jcyuan add  
                state <= STATE_IDLE;//jcyuan add
end

//---------------------------------------------
//------------Register transfers---------------
//---------------------------------------------

//-------------------for index----------------
always @ (posedge RST or negedge SCL)
begin
        if (RST)
                index_pointer <= 8'h00;
        else if (stop_detect)
                index_pointer <= 8'h00;
        else if (ack_bit)//at the 9th bit -ack, the input_shift has one bytes
        begin
                if (state == STATE_IDX_PTR) //at the state get the inner-register index
                        index_pointer <= input_shift;
                else//ready for next read/write;bulk transfer of a block of data 
                        index_pointer <= index_pointer + 8'h01;
        end
end

//----------------for write---------------------------
//we only define 4 registers for operation
always @ (posedge RST or negedge SCL)
begin
        if (RST)
        begin
                reg_00 <= 8'h00;
                reg_01 <= 8'h00;
                reg_02 <= 8'h00;
        end//the moment the input_shift has one byte=8bits
        else if (write_strobe && (index_pointer == 8'h00))
                reg_00 <= input_shift;
        else if (write_strobe && (index_pointer == 8'h01))
                reg_01 <= input_shift;
        else if (write_strobe && (index_pointer == 8'h02))
                reg_02 <= input_shift;

end
assign reg_sel_in = reg_00[1:0];
always@(*) begin 
    if(reg_sel_in == 2'b00) begin
        conv = {reg_01,reg_02};
    end
    if(reg_sel_in == 2'b01) begin
        conf = {reg_01,reg_02};
    end
    if(reg_sel_in == 2'b10) begin
        lot = {reg_01,reg_02};
    end
    if(reg_sel_in == 2'b11) begin
        hit = {reg_01,reg_02};
    end
end
 

//------------------------for read-----------------------

assign sel = conf[14:12];

always @(*) begin
    conv_loaded = 0; // default
    if      (sel == 3'd0) begin conv[15:4] = i1; conv_loaded = 1; end
    else if (sel == 3'd1) begin conv[15:4] = i2; conv_loaded = 1; end
    else if (sel == 3'd2) begin conv[15:4] = i3; conv_loaded = 1; end
    else if (sel == 3'd3) begin conv[15:4] = i4; conv_loaded = 1; end
    else if (sel == 3'd4) begin conv[15:4] = i5; conv_loaded = 1; end
    else if (sel == 3'd5) begin conv[15:4] = i6; conv_loaded = 1; end
    else if (sel == 3'd6) begin conv[15:4] = i7; conv_loaded = 1; end
    else if (sel == 3'd7) begin conv[15:4] = i8; conv_loaded = 1; end
    else                  begin conv[15:4] = 12'd0; conv_loaded = 0; end
end


assign reg_sel_in = reg_00[1:0];
always@(*) begin 
    if(reg_sel_in == 2'b00) begin
        reg_01 = conv[15:8];
        reg_02 = conv[7:0];
    end
    if(reg_sel_in == 2'b01) begin
        reg_01 = conf[15:8];
        reg_02 = conf[7:0];
    end
    if(reg_sel_in == 2'b10) begin
        reg_01 = lot[15:8];
        reg_02 = lot[7:0];
    end
    if(reg_sel_in == 2'b11) begin
        reg_01 = hit[15:8];
        reg_02 = hit[7:0];
    end
end

always @ (negedge SCL)
begin   
        if (lsb_bit)//at one byte that can be load the output_shift
        begin   
                case (index_pointer)
                8'h00: output_shift <= reg_01;
                8'h01: output_shift <= reg_02;
                
                endcase
        end
        else
                output_shift <= {output_shift[6:0], 1'b0};
                //once the shift it,after 8 times the output_shift=8'b0
                //the 9th bit is 0 for the RESTART for address match slave ACK 
end

//---------------------------------------------
//------------Output driver--------------------
//---------------------------------------------

always @ (posedge RST or negedge SCL)
begin   
        if (RST)
                output_control <= 1'b1;
        else if (start_detect)
                output_control <= 1'b1;
        else if (lsb_bit)
        begin   
                output_control <=
                    !(((state == STATE_DEV_ADDR) && address_detect) ||
                      (state == STATE_IDX_PTR) ||
                      (state == STATE_WRITE)); 
                //when operation is wirte 
                //addr match gen ACK,the index get gen ACK,and write data gen ACK
        end
        else if (ack_bit)
        begin
                // Deliver the first bit of the next slave-to-master
                // transfer, if applicable.
                if (((state == STATE_READ) && master_ack) ||
                    ((state == STATE_DEV_ADDR) &&
                        address_detect && read_write_bit))
                        output_control <= output_shift[7];
                        //for the RESTART and send the addr ACK for 1'b0
                        //for the read and master ack both slave is pull down
                else
                        output_control <= 1'b1;
        end
        else if (state == STATE_READ)//for read send output shift to SDA
                output_control <= output_shift[7];
        else
                output_control <= 1'b1;
end
endmodule